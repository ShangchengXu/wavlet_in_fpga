module wavlet(
	input clk,
	input rst_n,
	input [15:0] data_in,
	output [19:0] data_out
)