interface wavlet_interface_inner;




endinterface