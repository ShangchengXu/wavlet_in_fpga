interface wavlet_interface_port;
logic clk;
logic rst_n;
logic [15:0] data_in;
logic [20:0] data_out_hd;
logic [20:0] data_out_ld;




endinterface